`timescale 1ns / 1ps

module debounce(
    input clk,          // 100MHz clock
    input btn_in,       // ��������ԧ
    output reg btn_out  // �ѭ�ҳ����ͧ���� (Pulse 1 ����)
    );

    reg [19:0] count;
    reg btn_prev;
    reg btn_stable;

    always @(posedge clk) begin
        // ����ѭ�ҳ����¹ ���������Ѻ����
        if (btn_in != btn_stable) begin
            count <= count + 1;
            // ��ҹ�觹ҹ�� (����ҳ 10ms) �������Ѻ�������
            if (count == 20'd1_000_000) begin
                btn_stable <= btn_in;
                count <= 0;
            end
        end else begin
            count <= 0;
        end
        
        // ���ҧ�ѭ�ҳ Pulse ��§ 1 clock cycle ����͡�����
        btn_prev <= btn_stable;
        btn_out <= (btn_stable == 1'b1 && btn_prev == 1'b0) ? 1'b1 : 1'b0;
    end
endmodule