`timescale 1ns / 1ps
module top(
    input clk,          // Clock 100MHz
    input btnC,         // ������ҧ = ���ⴴ (Jump)
    input btnL,         // [NEW] �������� = �������/��ʵ��� (Start)
    input sw0,          // ��Ե�� 0 = ���絺��� (Reset)
    output [3:0] vgaRed,
    output [3:0] vgaGreen,
    output [3:0] vgaBlue,
    output Hsync,
    output Vsync,
    output [6:0] seg,   // 7-segment cathodes
    output [3:0] an     // 7-segment anodes
    );

    wire clean_jump;    // �ѭ�ҳ���ⴴ��� Debounce ����
    wire clean_start;   // [NEW] �ѭ�ҳ���������� Debounce ����
    
    wire video_on;
    wire [9:0] x, y;
    wire [11:0] rgb_out;
    wire [13:0] score;
    wire p_tick;

    // 1. Instantiate Debouncers
    // ��Ƿ�� 1: ����Ѻ�������ⴴ (btnC)
    debounce db_jump (
        .clk(clk),
        .btn_in(btnC),
        .btn_out(clean_jump)
    );
    
    // [NEW] ��Ƿ�� 2: ����Ѻ����������� (btnL)
    debounce db_start (
        .clk(clk),
        .btn_in(btnL),
        .btn_out(clean_start)
    );

    // 2. Instantiate VGA Controller
    vga_display vga_inst (
        .clk(clk),
        .rst(sw0),
        .hsync(Hsync),
        .vsync(Vsync),
        .video_on(video_on),
        .x(x),
        .y(y),
        .p_tick(p_tick)
    );

    // 3. Instantiate Game Engine
    game_engine game_inst (
        .clk(clk),          
        .rst(sw0),
        .jump_btn(clean_jump),   // ������������ⴴ
        .start_btn(clean_start), // [NEW] ����������������
        .video_on(video_on),
        .pixel_x(x),
        .pixel_y(y),
        .rgb(rgb_out),
        .score(score)
    );

    // 4. Instantiate 7-Segment Display
    seg7_control seg_inst (
        .clk(clk),
        .number(score),
        .an(an),
        .seg(seg)
    );

    // ������ѭ�ҳ���͡ VGA Port
    assign vgaRed   = rgb_out[11:8];
    assign vgaGreen = rgb_out[7:4];
    assign vgaBlue  = rgb_out[3:0];

endmodule