`timescale 1ns / 1ps

module vga_tb;

    // ==========================================
    // 1. ��С�ȵ����
    // ==========================================
    reg clk;
    reg rst;

    // Outputs �ҡ Module VGA
    wire hsync;
    wire vsync;
    wire video_on;
    wire [9:0] x;
    wire [9:0] y;
    wire p_tick;

    // ==========================================
    // 2. �������͡Ѻ vga_display (Instantiate)
    // ==========================================
    vga_display uut (
        .clk(clk),
        .rst(rst),
        .hsync(hsync),
        .vsync(vsync),
        .video_on(video_on),
        .x(x),
        .y(y),
        .p_tick(p_tick)
    );

    // ==========================================
    // 3. ���ҧ Clock 100MHz (�Ӥѭ�ҡ!)
    // ==========================================
    initial begin
        clk = 0;
        // ��Ѻ��ҷء 5ns -> �Һ 10ns -> 100MHz
        forever #5 clk = ~clk; 
    end

    // ==========================================
    // 4. ��ǹ��Ǩ�ͺ�� (Monitor) [NEW!]
    // ==========================================
    // ��ǹ���Ъ��¾�����ͤ����͡������� V-Sync ��ŧ��
    initial begin
        // �����鹪�ǧ Reset ��͹
        #200; 
        
        // ǹ�ٻ�ͨѺ�ѭ�ҳ V-Sync ��ŧ (negedge)
        forever begin
            @(negedge vsync); 
            $display("Time: %t | V-Sync Detected! (Frame End)", $time);
        end
    end

    // ==========================================
    // 5. �ӴѺ��÷��ͺ (Stimulus)
    // ==========================================
    initial begin
        // �������: ��駤��������� ��С� Reset
        $display("Simulation Start...");
        rst = 1; 
        
        // �� 100ns ���ǻ���� Reset
        #100;
        rst = 0;
        $display("Reset Released. VGA Running...");

        // �ѹ���� ����ҳ 35ms (���������� V-Sync ���ҧ���� 2 �ͺ)
        // 1 ms = 1,000,000 ns
        #35000000; 

        $display("Simulation Timeout. Finishing...");
        $finish;
    end

endmodule